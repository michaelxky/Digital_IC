* SPICE NETLIST
***************************************

.SUBCKT GREYCELLHP Ph Gl Gh VDD GND GG
** N=9 EP=6 IP=0 FDC=8
M0 9 Ph GND GND NMOS_VTG L=5e-08 W=9e-08 AD=1.7775e-14 AS=1.1475e-14 PD=5.75e-07 PS=4.35e-07 $X=2490 $Y=2135 $D=5
M1 5 Gl 9 GND NMOS_VTG L=5e-08 W=9e-08 AD=2.3175e-14 AS=1.7775e-14 PD=6.95e-07 PS=5.75e-07 $X=2985 $Y=2135 $D=5
M2 GND Gh 5 GND NMOS_VTG L=5e-08 W=9e-08 AD=1.2825e-14 AS=2.3175e-14 PD=4.65e-07 PS=6.95e-07 $X=3600 $Y=2135 $D=5
M3 GG 5 GND GND NMOS_VTG L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=4355 $Y=2135 $D=5
M4 VDD Ph 3 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=3.555e-14 AS=2.25e-14 PD=7.55e-07 PS=6.1e-07 $X=2490 $Y=3115 $D=4
M5 3 Gl VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=4.635e-14 AS=3.555e-14 PD=8.75e-07 PS=7.55e-07 $X=2985 $Y=3115 $D=4
M6 5 Gh 3 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=2.565e-14 AS=4.635e-14 PD=6.45e-07 PS=8.75e-07 $X=3600 $Y=3115 $D=4
M7 GG 5 VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=4355 $Y=3115 $D=4
.ENDS
***************************************
