* SPICE NETLIST
***************************************

.SUBCKT BLACK Pl Ph Pout Gl Gh Gout VDD GND
** N=13 EP=8 IP=0 FDC=14
M0 12 Pl GND GND NMOS_VTG L=5e-08 W=9e-08 AD=1.305e-14 AS=9.45e-15 PD=4.7e-07 PS=3.9e-07 $X=360 $Y=560 $D=5
M1 2 Ph 12 GND NMOS_VTG L=5e-08 W=9e-08 AD=9.45e-15 AS=1.305e-14 PD=3.9e-07 PS=4.7e-07 $X=750 $Y=560 $D=5
M2 Pout 2 GND GND NMOS_VTG L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=1510 $Y=560 $D=5
M3 13 Ph GND GND NMOS_VTG L=5e-08 W=9e-08 AD=1.7775e-14 AS=1.1475e-14 PD=5.75e-07 PS=4.35e-07 $X=2320 $Y=535 $D=5
M4 9 Gl 13 GND NMOS_VTG L=5e-08 W=9e-08 AD=2.61e-14 AS=1.7775e-14 PD=7.6e-07 PS=5.75e-07 $X=2815 $Y=535 $D=5
M5 GND Gh 9 GND NMOS_VTG L=5e-08 W=9e-08 AD=1.2825e-14 AS=2.61e-14 PD=4.65e-07 PS=7.6e-07 $X=3495 $Y=535 $D=5
M6 Gout 9 GND GND NMOS_VTG L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=4290 $Y=560 $D=5
M7 2 Pl VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=2.61e-14 AS=1.89e-14 PD=6.5e-07 PS=5.7e-07 $X=360 $Y=1540 $D=4
M8 VDD Ph 2 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.61e-14 PD=5.7e-07 PS=6.5e-07 $X=750 $Y=1540 $D=4
M9 Pout 2 VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=1510 $Y=1540 $D=4
M10 VDD Ph 8 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=3.555e-14 AS=2.25e-14 PD=7.55e-07 PS=6.1e-07 $X=2320 $Y=1515 $D=4
M11 8 Gl VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=5.22e-14 AS=3.555e-14 PD=9.4e-07 PS=7.55e-07 $X=2815 $Y=1515 $D=4
M12 9 Gh 8 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=2.475e-14 AS=5.22e-14 PD=6.35e-07 PS=9.4e-07 $X=3495 $Y=1515 $D=4
M13 Gout 9 VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=4290 $Y=1540 $D=4
.ENDS
***************************************
