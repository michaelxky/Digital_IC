* SPICE NETLIST
***************************************

.SUBCKT AOI21 B OUT A2 VDD A1 GND
** N=8 EP=6 IP=0 FDC=6
M0 OUT B GND GND NMOS_VTG L=5e-08 W=9e-08 AD=2.61e-14 AS=1.2825e-14 PD=7.6e-07 PS=4.65e-07 $X=400 $Y=640 $D=5
M1 8 A2 OUT GND NMOS_VTG L=5e-08 W=9e-08 AD=1.7775e-14 AS=2.61e-14 PD=5.75e-07 PS=7.6e-07 $X=1080 $Y=640 $D=5
M2 GND A1 8 GND NMOS_VTG L=5e-08 W=9e-08 AD=1.1475e-14 AS=1.7775e-14 PD=4.35e-07 PS=5.75e-07 $X=1575 $Y=640 $D=5
M3 6 B OUT VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=5.22e-14 AS=2.475e-14 PD=9.4e-07 PS=6.35e-07 $X=400 $Y=1620 $D=4
M4 VDD A2 6 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=3.555e-14 AS=5.22e-14 PD=7.55e-07 PS=9.4e-07 $X=1080 $Y=1620 $D=4
M5 6 A1 VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=2.25e-14 AS=3.555e-14 PD=6.1e-07 PS=7.55e-07 $X=1575 $Y=1620 $D=4
.ENDS
***************************************
