* SPICE NETLIST
***************************************

.SUBCKT INVX2 IN OUT GND VDD
** N=4 EP=4 IP=0 FDC=4
M0 OUT IN GND GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=355 $Y=490 $D=5
M1 GND IN OUT GND NMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=735 $Y=490 $D=5
M2 OUT IN VDD VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.2e-14 AS=3.45e-14 PD=8.8e-07 PS=8.3e-07 $X=355 $Y=1280 $D=4
M3 VDD IN OUT VDD PMOS_VTG L=5e-08 W=3e-07 AD=3.15e-14 AS=4.2e-14 PD=8.1e-07 PS=8.8e-07 $X=735 $Y=1280 $D=4
.ENDS
***************************************
