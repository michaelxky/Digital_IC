* SPICE NETLIST
***************************************

.SUBCKT AND B A VDD GND OUT
** N=7 EP=5 IP=0 FDC=6
M0 7 B GND GND NMOS_VTG L=5e-08 W=9e-08 AD=1.305e-14 AS=9.45e-15 PD=4.7e-07 PS=3.9e-07 $X=360 $Y=520 $D=5
M1 1 A 7 GND NMOS_VTG L=5e-08 W=9e-08 AD=9.45e-15 AS=1.305e-14 PD=3.9e-07 PS=4.7e-07 $X=750 $Y=520 $D=5
M2 OUT 1 GND GND NMOS_VTG L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=1510 $Y=520 $D=5
M3 1 B VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=2.61e-14 AS=1.89e-14 PD=6.5e-07 PS=5.7e-07 $X=360 $Y=1500 $D=4
M4 VDD A 1 VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.61e-14 PD=5.7e-07 PS=6.5e-07 $X=750 $Y=1500 $D=4
M5 OUT 1 VDD VDD PMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=1510 $Y=1500 $D=4
.ENDS
***************************************
