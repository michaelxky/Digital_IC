* SPICE NETLIST
***************************************

.SUBCKT DBUFFER IN OUT GND VDD
** N=5 EP=4 IP=0 FDC=16
M0 2 IN GND GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.07e-14 PD=6.4e-07 PS=5.9e-07 $X=2045 $Y=1030 $D=5
M1 GND IN 2 GND NMOS_VTG L=5e-08 W=1.8e-07 AD=3.465e-14 AS=2.52e-14 PD=7.45e-07 PS=6.4e-07 $X=2425 $Y=1030 $D=5
M2 OUT 2 GND GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.52e-14 AS=3.465e-14 PD=6.4e-07 PS=7.45e-07 $X=2910 $Y=1030 $D=5
M3 GND 2 OUT GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.7e-14 AS=2.52e-14 PD=6.6e-07 PS=6.4e-07 $X=3290 $Y=1030 $D=5
M4 OUT 2 GND GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.7e-14 PD=6.4e-07 PS=6.6e-07 $X=3690 $Y=1030 $D=5
M5 GND 2 OUT GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.52e-14 PD=6.8e-07 PS=6.4e-07 $X=4070 $Y=1030 $D=5
M6 OUT 2 GND GND NMOS_VTG L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.88e-14 PD=6.4e-07 PS=6.8e-07 $X=4490 $Y=1030 $D=5
M7 GND 2 OUT GND NMOS_VTG L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=4870 $Y=1030 $D=5
M8 2 IN VDD VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.2e-14 AS=3.45e-14 PD=8.8e-07 PS=8.3e-07 $X=2045 $Y=1820 $D=4
M9 VDD IN 2 VDD PMOS_VTG L=5e-08 W=3e-07 AD=5.775e-14 AS=4.2e-14 PD=9.85e-07 PS=8.8e-07 $X=2425 $Y=1820 $D=4
M10 OUT 2 VDD VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.2e-14 AS=5.775e-14 PD=8.8e-07 PS=9.85e-07 $X=2910 $Y=1820 $D=4
M11 VDD 2 OUT VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.5e-14 AS=4.2e-14 PD=9e-07 PS=8.8e-07 $X=3290 $Y=1820 $D=4
M12 OUT 2 VDD VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.2e-14 AS=4.5e-14 PD=8.8e-07 PS=9e-07 $X=3690 $Y=1820 $D=4
M13 VDD 2 OUT VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.8e-14 AS=4.2e-14 PD=9.2e-07 PS=8.8e-07 $X=4070 $Y=1820 $D=4
M14 OUT 2 VDD VDD PMOS_VTG L=5e-08 W=3e-07 AD=4.2e-14 AS=4.8e-14 PD=8.8e-07 PS=9.2e-07 $X=4490 $Y=1820 $D=4
M15 VDD 2 OUT VDD PMOS_VTG L=5e-08 W=3e-07 AD=3.15e-14 AS=4.2e-14 PD=8.1e-07 PS=8.8e-07 $X=4870 $Y=1820 $D=4
.ENDS
***************************************
